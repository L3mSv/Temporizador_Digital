library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity display24 is
  port (
  ) ;
end display24; 

architecture arq of display24 is

begin

end arq ;